* EESchema Netlist Version 1.1 (Spice format) creation date: 07/05/2014 10:33:00

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
V1  ? ? VSOURCE		
R1  ? ? R		

.end
